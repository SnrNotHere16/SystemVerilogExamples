`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// File:AssertionsPracticeTB2.sv
// output 
//init time start: 0

//Time: 5 ns Started: 5 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 15 ns Started: 15 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 25 ns Started: 25 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 35 ns Started: 35 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 45 ns Started: 45 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 55 ns Started: 55 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 65 ns Started: 65 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 75 ns Started: 75 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 85 ns Started: 85 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 95 ns Started: 95 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 105 ns Started: 105 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 115 ns Started: 115 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 125 ns Started: 125 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 135 ns Started: 135 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 145 ns Started: 145 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Trigger pass time start: 150.00 ns

//Time: 155 ns Started: 155 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 165 ns Started: 165 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 175 ns Started: 175 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 185 ns Started: 185 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 195 ns Started: 165 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:1 b:1

//Time: 195 ns Started: 195 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 205 ns Started: 175 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:1 b:1

//Time: 205 ns Started: 205 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 215 ns Started: 185 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 215 ns Started: 215 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 225 ns Started: 195 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 225 ns Started: 225 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 235 ns Started: 205 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 235 ns Started: 235 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 245 ns Started: 245 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 255 ns Started: 255 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 265 ns Started: 265 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Trigger fail time start: 270.00 ns

//Time: 275 ns Started: 275 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 285 ns Started: 285 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 295 ns Started: 285 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b failed: a:1 b:0

//Time: 295 ns Started: 295 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 305 ns Started: 295 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b failed: a:1 b:0

//Time: 305 ns Started: 305 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 315 ns Started: 305 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b failed: a:1 b:0

//Time: 315 ns Started: 315 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 325 ns Started: 325 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 335 ns Started: 335 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 345 ns Started: 315 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 345 ns Started: 345 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 355 ns Started: 325 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 355 ns Started: 355 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 365 ns Started: 335 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:72
//a_b passed: a:0 b:1

//Time: 365 ns Started: 365 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Use not pass start time: 370.00 ns

//Time: 375 ns Started: 375 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:x d:x

//Time: 385 ns Started: 385 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:0 d:0

//Time: 395 ns Started: 395 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:0 d:0

//Time: 405 ns Started: 405 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:0 d:0

//Time: 415 ns Started: 415 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:0 d:0

//Time: 435 ns Started: 425 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:1 d:0

//Use not fail start time1: 440.00 ns

//Time: 445 ns Started: 435 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:1 d:0

//Time: 455 ns Started: 445 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d failed: c:1 d:1

//Time: 465 ns Started: 455 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d failed: c:1 d:1

//Time: 475 ns Started: 465 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d failed: c:1 d:1

//Use not fail start time2: 480.00 ns

//Time: 485 ns Started: 475 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d failed: c:1 d:1

//Time: 495 ns Started: 485 ns Scope: /AssertionsPracticeTB2 File: /home/user/Desktop/VivadoEX/Sample/Sample.srcs/sources_1/new/AssertionsPracticeTB2.sv Line:73
//c_d passed: c:1 d:0
//$stop called at time : 500 ns
//////////////////////////////////////////////////////////////////////////////////


module AssertionsPracticeTB2();
    logic clk, reset; 
    logic a,b,c,d,e,f,g; 
     
    task init(); 
        $display ("\ninit time start: %0t", $realtime);
        repeat (10) @ (negedge clk) begin reset <= 1'b1; a <= 1; b <= 0;  end
        repeat (5) @ (negedge clk) begin reset <= 1'b0; a <= 0; b <= 0; end 
    endtask: init
    
    initial begin 
        clk = 1'b0; 
    end 

    always#5 clk = ~clk; 
    
    initial begin 
        init(); 
        // trigger pass 
        $timeformat(-9, 2, " ns", 20);
        $display ("\nTrigger pass time start: %0t", $realtime);
        repeat (5) @ (negedge clk) begin a <= 1; b <= 1; end 
        repeat (5) @ (negedge clk) begin a <= 0; b <= 1; end 
        repeat (2) @ (negedge clk) begin a <= 0; b <= 0; end 
        
        //trigger fail 
        $display ("\nTrigger fail time start: %0t", $realtime);
        repeat (4) @ (negedge clk) begin a <= 1; b <= 0; end 
        repeat (2) @ (negedge clk) begin  b <= 1; end 
        repeat (4) @ (negedge clk) begin a <= 0; end 
        
        //Use not pass 
        $display ("\nUse not pass start time: %0t", $realtime);
        repeat (4) @ (negedge clk) begin c <= 0; d <= 0; end 
        repeat (3) @ (negedge clk) begin c <= 1; d <= 0; end 
        
        //Use not fail 
        $display ("\nUse not fail start time1: %0t", $realtime);
        repeat (4) @ (negedge clk) begin c <= 1; d <= 1; end 
        $display ("\nUse not fail start time2: %0t", $realtime);
        repeat (2) @ (negedge clk) d <= 0; 
        $stop; 
    end    
   
   
   sequence a_b_s; 
//        ## 1 b == 0 ## 1 b == 0 ## 1 b == 0 ## 1 b == 0;
          ##1 b[*3]; 
//        ##1 b[->3]; //go to repetition 
//        ##1 b[=3]; //non-consecutive repetition 
   endsequence: a_b_s 
   
   property a_b_p; 
         @ (posedge clk) disable iff (reset) a |-> a_b_s; 
   endproperty: a_b_p
   
 sequence c_d_s;
    @ (posedge clk) c ##1 d;
 endsequence: c_d_s
 
 property c_d_p;
    not c_d_s; 
 endproperty: c_d_p
 
   a_b_ap:assert property (a_b_p) $display ("a_b passed: a:%d b:%d", a, b); else $display ("a_b failed: a:%d b:%d", a, b); 
   c_d_ap: assert property (c_d_p) $display ("c_d passed: c:%d d:%d", c, d); else $display ("c_d failed: c:%d d:%d", c, d);
endmodule
