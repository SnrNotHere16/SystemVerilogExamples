`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// File: FunctionalCoverageTB3.sv
// output: 

//# coverPClass created
//# 
//# Begin
//# ** Note: $stop    : testbench.sv(46)
//#    Time: 125 ns  Iteration: 1  Instance: /FunctionalCoverageTB7
//# Break in Module FunctionalCoverageTB7 at testbench.sv line 46
//# Coverage Report by instance with details
//# 
//# =================================================================================
//# === Instance: /FunctionalCoverageTB7
//# === Design Unit: work.FunctionalCoverageTB7
//# =================================================================================
//# 
//# Covergroup Coverage:
//#     Covergroups                      2        na        na    10.00%
//#         Coverpoints/Crosses          4        na        na        na
//#             Covergroup Bins         42         4        38     9.52%
//# ----------------------------------------------------------------------------------------------------------
//# Covergroup                                             Metric       Goal       Bins    Status               
//#                                                                                                          
//# ----------------------------------------------------------------------------------------------------------
//#  TYPE /FunctionalCoverageTB7/coverPClass/a_c           20.00%        100          -    Uncovered            
//#     covered/total bins:                                     4         18          -                      
//#     missing/total bins:                                    14         18          -                      
//#     % Hit:                                             22.22%        100          -                      
//#     Coverpoint a1                                      40.00%        100          -    Uncovered            
//#         covered/total bins:                                 4         10          -                      
//#         missing/total bins:                                 6         10          -                      
//#         % Hit:                                         40.00%        100          -                      
//#     Coverpoint c1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#  Covergroup instance \/FunctionalCoverageTB7/coverPClass::a_c  
//#                                                        20.00%        100          -    Uncovered            
//#     covered/total bins:                                     4         18          -                      
//#     missing/total bins:                                    14         18          -                      
//#     % Hit:                                             22.22%        100          -                      
//#     Coverpoint a1                                      40.00%        100          -    Uncovered            
//#         covered/total bins:                                 4         10          -                      
//#         missing/total bins:                                 6         10          -                      
//#         % Hit:                                         40.00%        100          -                      
//#         bin a0[0]                                           0          1          -    ZERO                 
//#         bin a0[3]                                           4          1          -    Covered              
//#         bin a0[6]                                           1          1          -    Covered              
//#         bin a0[9]                                           0          1          -    ZERO                 
//#         bin at0                                             2          1          -    Covered              
//#         bin at1                                             0          1          -    ZERO                 
//#         bin at2                                             4          1          -    Covered              
//#         bin at3                                             0          1          -    ZERO                 
//#         bin at4                                             0          1          -    ZERO                 
//#         bin at5                                             0          1          -    ZERO                 
//#     Coverpoint c1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//#  TYPE /FunctionalCoverageTB7/coverPClass/b_e_d          0.00%        100          -    ZERO                 
//#     covered/total bins:                                     0         24          -                      
//#     missing/total bins:                                    24         24          -                      
//#     % Hit:                                              0.00%        100          -                      
//#     Coverpoint b1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0         16          -                      
//#         missing/total bins:                                16         16          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//#         bin auto[8]                                         0          1          -    ZERO                 
//#         bin auto[9]                                         0          1          -    ZERO                 
//#         bin auto[10]                                        0          1          -    ZERO                 
//#         bin auto[11]                                        0          1          -    ZERO                 
//#         bin auto[12]                                        0          1          -    ZERO                 
//#         bin auto[13]                                        0          1          -    ZERO                 
//#         bin auto[14]                                        0          1          -    ZERO                 
//#         bin auto[15]                                        0          1          -    ZERO                 
//#     Coverpoint dPe                                      0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//# 
//# COVERGROUP COVERAGE:
//# ----------------------------------------------------------------------------------------------------------
//# Covergroup                                             Metric       Goal       Bins    Status               
//#                                                                                                          
//# ----------------------------------------------------------------------------------------------------------
//#  TYPE /FunctionalCoverageTB7/coverPClass/a_c           20.00%        100          -    Uncovered            
//#     covered/total bins:                                     4         18          -                      
//#     missing/total bins:                                    14         18          -                      
//#     % Hit:                                             22.22%        100          -                      
//#     Coverpoint a1                                      40.00%        100          -    Uncovered            
//#         covered/total bins:                                 4         10          -                      
//#         missing/total bins:                                 6         10          -                      
//#         % Hit:                                         40.00%        100          -                      
//#     Coverpoint c1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#  Covergroup instance \/FunctionalCoverageTB7/coverPClass::a_c  
//#                                                        20.00%        100          -    Uncovered            
//#     covered/total bins:                                     4         18          -                      
//#     missing/total bins:                                    14         18          -                      
//#     % Hit:                                             22.22%        100          -                      
//#     Coverpoint a1                                      40.00%        100          -    Uncovered            
//#         covered/total bins:                                 4         10          -                      
//#         missing/total bins:                                 6         10          -                      
//#         % Hit:                                         40.00%        100          -                      
//#         bin a0[0]                                           0          1          -    ZERO                 
//#         bin a0[3]                                           4          1          -    Covered              
//#         bin a0[6]                                           1          1          -    Covered              
//#         bin a0[9]                                           0          1          -    ZERO                 
//#         bin at0                                             2          1          -    Covered              
//#         bin at1                                             0          1          -    ZERO                 
//#         bin at2                                             4          1          -    Covered              
//#         bin at3                                             0          1          -    ZERO                 
//#         bin at4                                             0          1          -    ZERO                 
//#         bin at5                                             0          1          -    ZERO                 
//#     Coverpoint c1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//#  TYPE /FunctionalCoverageTB7/coverPClass/b_e_d          0.00%        100          -    ZERO                 
//#     covered/total bins:                                     0         24          -                      
//#     missing/total bins:                                    24         24          -                      
//#     % Hit:                                              0.00%        100          -                      
//#     Coverpoint b1                                       0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0         16          -                      
//#         missing/total bins:                                16         16          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//#         bin auto[8]                                         0          1          -    ZERO                 
//#         bin auto[9]                                         0          1          -    ZERO                 
//#         bin auto[10]                                        0          1          -    ZERO                 
//#         bin auto[11]                                        0          1          -    ZERO                 
//#         bin auto[12]                                        0          1          -    ZERO                 
//#         bin auto[13]                                        0          1          -    ZERO                 
//#         bin auto[14]                                        0          1          -    ZERO                 
//#         bin auto[15]                                        0          1          -    ZERO                 
//#     Coverpoint dPe                                      0.00%        100          -    ZERO                 
//#         covered/total bins:                                 0          8          -                      
//#         missing/total bins:                                 8          8          -                      
//#         % Hit:                                          0.00%        100          -                      
//#         bin auto[0]                                         0          1          -    ZERO                 
//#         bin auto[1]                                         0          1          -    ZERO                 
//#         bin auto[2]                                         0          1          -    ZERO                 
//#         bin auto[3]                                         0          1          -    ZERO                 
//#         bin auto[4]                                         0          1          -    ZERO                 
//#         bin auto[5]                                         0          1          -    ZERO                 
//#         bin auto[6]                                         0          1          -    ZERO                 
//#         bin auto[7]                                         0          1          -    ZERO                 
//# 
//# TOTAL COVERGROUP COVERAGE: 10.00%  COVERGROUP TYPES: 2
//# 
//# Total Coverage By Instance (filtered view): 10.00%
//////////////////////////////////////////////////////////////////////////////////


module FunctionalCoverageTB7(); 
	logic clk; 
  	logic rest; 
  	logic reset; 
	class coverPClass; 
	  logic [3:0] a,b; 
      logic [2:0] c, d, e, f; 
		covergroup a_c @(posedge clk);  
          a1: coverpoint a {
            bins a0 [] = {[0:10]} with (item%3 == 0); //divides the bins into only values that fufill the statement, 4 bins
            bins at0 = (3[*3]); // 3=>3=>3, 3 consecutive 3s 
            bins at1 = (4[*3:5]); //( 4=>4=>4 ), ( 4=>4=>4=>4 ), ( 4=>4=>4=>4=>4 ) 3  to 5 consecutive 4s 
            bins at2 = (5 [= 2]);//nonconsecutive 2 5's 
            bins at3 = (4 => 5 => 6), ([7:9],10=>11,12); // 4=>5=>6, or 7=>11, 8=>11, 9=>11, 10=>11, 7=>12, 8=>12, 9=>12, 10=>12.
            bins at4 = (12 => 3 [-> 1]); // 12 => ....3 nonconsecutive 3 
            bins at5 = ( 2 [-> 3:5] );// 3 to 5 nonconsectuive 2s 
          } 
          c1: coverpoint c; 
          	//aXc: cross a,c; 
        endgroup: a_c
		
      covergroup b_e_d; 
        	b1: coverpoint b iff (!reset);
        	dPe: coverpoint d+e; 
		endgroup: b_e_d
		
		function new(); 
			$display("coverPClass created\n");
			a_c = new(); 
            b_e_d = new(); 
		endfunction: new 
	endclass: coverPClass 
	
  	initial begin 
    	clk = 1'b0; 
    end 
	always #5 clk = ~clk; 
  	coverPClass cov = new(); 
	initial begin 
      $display("Begin");  
      repeat (4) @(posedge clk) cov.a <= 3;  
      @ (posedge clk) cov.a <= 5; 
      repeat(3) @ (posedge clk) cov.a <= cov.a+1; 
      repeat (2) @(posedge clk) cov.a <= 5; 

      $stop; 
    end 
  
  

endmodule: FunctionalCoverageTB7 