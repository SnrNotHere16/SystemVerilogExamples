module FunctionalCoverageTB5();
	



endmodule: FunctionalCoverageTB5