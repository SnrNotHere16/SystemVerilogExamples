module FunctionalCoverageTB7(); 






endmodule: FunctionalCoverageTB7 