//////////////////////////////////////////////////////////////////////////////////
// File: FunctionalCoverageTB4.sv
// Output: 
// # do run.do
//# Begin
//# Coverage Report by instance with details
//# 
//# =================================================================================
//# === Instance: /FunctionalCoverageTB4
//# === Design Unit: work.FunctionalCoverageTB4
//# =================================================================================
//# 
//# Covergroup Coverage:
//#     Covergroups                      1        na        na    73.07%
//#         Coverpoints/Crosses          2        na        na        na
//#             Covergroup Bins         17        10         7    58.82%
//# ----------------------------------------------------------------------------------------------------------
//# Covergroup                                             Metric       Goal       Bins    Status               
//#                                                                                                          
//# ----------------------------------------------------------------------------------------------------------
//#  TYPE /FunctionalCoverageTB4/a_c                       73.07%        100          -    Uncovered            
//#     covered/total bins:                                    10         17          -                      
//#     missing/total bins:                                     7         17          -                      
//#     % Hit:                                             58.82%        100          -                      
//#     Coverpoint a_1                                     46.15%        100          -    Uncovered            
//#         covered/total bins:                                 6         13          -                      
//#         missing/total bins:                                 7         13          -                      
//#         % Hit:                                         46.15%        100          -                      
//#     Coverpoint c_1                                    100.00%        100          -    Covered              
//#         covered/total bins:                                 4          4          -                      
//#         missing/total bins:                                 0          4          -                      
//#         % Hit:                                        100.00%        100          -                      
//#  Covergroup instance \/FunctionalCoverageTB4/a_c_i  
//#                                                        73.07%        100          -    Uncovered            
//#     covered/total bins:                                    10         17          -                      
//#     missing/total bins:                                     7         17          -                      
//#     % Hit:                                             58.82%        100          -                      
//#     Coverpoint a_1                                     46.15%        100          -    Uncovered            
//#         covered/total bins:                                 6         13          -                      
//#         missing/total bins:                                 7         13          -                      
//#         % Hit:                                         46.15%        100          -                      
//#         bin a0                                              1          1          -    Covered              
//#         bin a1[0]                                           1          1          -    Covered              
//#         bin a1[1]                                           1          1          -    Covered              
//#         bin a1[2]                                           3          1          -    Covered              
//#         bin a2[8]                                           0          1          -    ZERO                 
//#         bin a2[9]                                           0          1          -    ZERO                 
//#         bin a2[10]                                          0          1          -    ZERO                 
//#         bin a2[11]                                          0          1          -    ZERO                 
//#         bin a2[12]                                          0          1          -    ZERO                 
//#         bin a2[13]                                          0          1          -    ZERO                 
//#         bin a2[14]                                          0          1          -    ZERO                 
//#         bin a3[0]                                           2          1          -    Covered              
//#         bin a3[1]                                           2          1          -    Covered              
//#         default bin a4                                      6                     -    Occurred             
//#     Coverpoint c_1                                    100.00%        100          -    Covered              
//#         covered/total bins:                                 4          4          -                      
//#         missing/total bins:                                 0          4          -                      
//#         % Hit:                                        100.00%        100          -                      
//#         bin c0                                              1          1          -    Covered              
//#         bin c1[0]                                           1          1          -    Covered              
//#         bin c1[1]                                           1          1          -    Covered              
//#         bin c1[2]                                           1          1          -    Covered              
//#         default bin c2                                     12                     -    Occurred             
//# 
//# COVERGROUP COVERAGE:
//# ----------------------------------------------------------------------------------------------------------
//# Covergroup                                             Metric       Goal       Bins    Status               
//#                                                                                                          
//# ----------------------------------------------------------------------------------------------------------
//#  TYPE /FunctionalCoverageTB4/a_c                       73.07%        100          -    Uncovered            
//#     covered/total bins:                                    10         17          -                      
//#     missing/total bins:                                     7         17          -                      
//#     % Hit:                                             58.82%        100          -                      
//#     Coverpoint a_1                                     46.15%        100          -    Uncovered            
//#         covered/total bins:                                 6         13          -                      
//#         missing/total bins:                                 7         13          -                      
//#         % Hit:                                         46.15%        100          -                      
//#     Coverpoint c_1                                    100.00%        100          -    Covered              
//#         covered/total bins:                                 4          4          -                      
//#         missing/total bins:                                 0          4          -                      
//#         % Hit:                                        100.00%        100          -                      
//#  Covergroup instance \/FunctionalCoverageTB4/a_c_i  
//#                                                        73.07%        100          -    Uncovered            
//#     covered/total bins:                                    10         17          -                      
//#     missing/total bins:                                     7         17          -                      
//#     % Hit:                                             58.82%        100          -                      
//#     Coverpoint a_1                                     46.15%        100          -    Uncovered            
//#         covered/total bins:                                 6         13          -                      
//#         missing/total bins:                                 7         13          -                      
//#         % Hit:                                         46.15%        100          -                      
//#         bin a0                                              1          1          -    Covered              
//#         bin a1[0]                                           1          1          -    Covered              
//#         bin a1[1]                                           1          1          -    Covered              
//#         bin a1[2]                                           3          1          -    Covered              
//#         bin a2[8]                                           0          1          -    ZERO                 
//#         bin a2[9]                                           0          1          -    ZERO                 
//#         bin a2[10]                                          0          1          -    ZERO                 
//#         bin a2[11]                                          0          1          -    ZERO                 
//#         bin a2[12]                                          0          1          -    ZERO                 
//#         bin a2[13]                                          0          1          -    ZERO                 
//#         bin a2[14]                                          0          1          -    ZERO                 
//#         bin a3[0]                                           2          1          -    Covered              
//#         bin a3[1]                                           2          1          -    Covered              
//#         default bin a4                                      6                     -    Occurred             
//#     Coverpoint c_1                                    100.00%        100          -    Covered              
//#         covered/total bins:                                 4          4          -                      
//#         missing/total bins:                                 0          4          -                      
//#         % Hit:                                        100.00%        100          -                      
//#         bin c0                                              1          1          -    Covered              
//#         bin c1[0]                                           1          1          -    Covered              
//#         bin c1[1]                                           1          1          -    Covered              
//#         bin c1[2]                                           1          1          -    Covered              
//#         default bin c2                                     12                     -    Occurred             
//# 
//# TOTAL COVERGROUP COVERAGE: 73.07%  COVERGROUP TYPES: 1
//# 
//# Total Coverage By Instance (filtered view): 73.07%
//////////////////////////////////////////////////////////////////////////////////

module FunctionalCoverageTB4();  
	logic [4:0] a,b; 
	logic [3:0] c,d; 
	logic [1:0] e,f; 

	covergroup a_c; 
		a_1: coverpoint a {
          	bins a0 = {0,1,2}; //a0 1 bin
          	bins a1 [3] = {3,4,[5:7]}; //a1 3 bins: {3,4, [5:7]}
          	bins a2 [] = {8,9, 10, [11:14]}; //a2 7 bins 
            bins a3 [2] = {[15:19]}; //a3 2 bins:  (15,16), (17,18,19)
			bins a4 = default; 
		} 
     	
      c_1: coverpoint c {
        bins c0 = {[0:5]};
        bins c1 [3] = {[9:13]};
        bins c2 = default; 
        
      } 
	endgroup: a_c
  
    task a_bins (); 
    	a = 0; 
        a_c_i.sample(); 
      	a = 3; 
        a_c_i.sample();
      repeat (4) begin 
        a++; 
        a_c_i.sample(); 
      end 
      //The default bins - a3[0] - 2, a3[1] - 2
      a = 15; 
      a_c_i.sample(); 
      a = 16; 
      a_c_i.sample(); 
	  a = 17; 
      a_c_i.sample(); 
	  a = 18; 
      a_c_i.sample(); 
      //The default bins - 2 
      a = 25; 
      a_c_i.sample(); 
      a_c_i.sample();
    endtask: a_bins  
  
 	task c_bins(); 
    	c = 0; 
      	a_c_i.sample();
      	c = 9; 
      	a_c_i.sample();
      	c = 10; 
        a_c_i.sample();
      	c = 11; 
        a_c_i.sample();
      	c = 6;
      	a_c_i.sample();
        c = 15; 
        a_c_i.sample();
    endtask: c_bins    
	a_c a_c_i = new(); 
	initial begin 
		$display("Begin"); 
      	a_bins; 
      	c_bins; 
	end 



endmodule: FunctionalCoverageTB4 